library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity end_screen is
  port(
		clk : in std_logic;
		y_in : in  unsigned(5 downto 0);
		x_in : in unsigned(6 downto 0);
		rgb : out std_logic_vector(5 downto 0)
  );
end end_screen;
architecture synth of end_screen is

signal addr: std_logic_vector(12 downto 0);

begin
		
addr <= std_logic_vector(y_in) & std_logic_vector(x_in);
process (clk)
begin
	if rising_edge(clk) then
			case addr is
                        when "0010100000011" => rgb <= "000000";
            when "0010100000100" => rgb <= "000000";
            when "0010100000101" => rgb <= "000000";
            when "0010100000110" => rgb <= "000000";
            when "0010100001101" => rgb <= "000000";
            when "0010100001110" => rgb <= "000000";
            when "0010100001111" => rgb <= "000000";
            when "0010100010000" => rgb <= "000000";
            when "0010100010101" => rgb <= "000000";
            when "0010100010110" => rgb <= "000000";
            when "0010100011011" => rgb <= "000000";
            when "0010100011100" => rgb <= "000000";
            when "0010100100001" => rgb <= "000000";
            when "0010100100010" => rgb <= "000000";
            when "0010100100011" => rgb <= "000000";
            when "0010100100100" => rgb <= "000000";
            when "0010100101001" => rgb <= "000000";
            when "0010100101010" => rgb <= "000000";
            when "0010100101011" => rgb <= "000000";
            when "0010100101100" => rgb <= "000000";
            when "0010100101101" => rgb <= "000000";
            when "0010100101110" => rgb <= "000000";
            when "0010100110101" => rgb <= "000000";
            when "0010100110110" => rgb <= "000000";
            when "0010100110111" => rgb <= "000000";
            when "0010100111000" => rgb <= "000000";
            when "0010100111101" => rgb <= "000000";
            when "0010100111110" => rgb <= "000000";
            when "0010100111111" => rgb <= "000000";
            when "0010101000000" => rgb <= "000000";
            when "0010101000001" => rgb <= "000000";
            when "0010101000010" => rgb <= "000000";
            when "0010101000011" => rgb <= "000000";
            when "0010101000100" => rgb <= "000000";
            when "0010101000101" => rgb <= "000000";
            when "0010101000110" => rgb <= "000000";
            when "0010101001010" => rgb <= "000000";
            when "0010101001011" => rgb <= "000000";
            when "0010101001100" => rgb <= "000000";
            when "0010101001101" => rgb <= "000000";
            when "0010101001110" => rgb <= "000000";
            when "0010110000011" => rgb <= "000000";
            when "0010110000100" => rgb <= "000000";
            when "0010110000101" => rgb <= "000000";
            when "0010110000110" => rgb <= "000000";
            when "0010110001101" => rgb <= "000000";
            when "0010110001110" => rgb <= "000000";
            when "0010110001111" => rgb <= "000000";
            when "0010110010000" => rgb <= "000000";
            when "0010110010101" => rgb <= "000000";
            when "0010110010110" => rgb <= "000000";
            when "0010110011011" => rgb <= "000000";
            when "0010110011100" => rgb <= "000000";
            when "0010110100001" => rgb <= "000000";
            when "0010110100010" => rgb <= "000000";
            when "0010110100011" => rgb <= "000000";
            when "0010110100100" => rgb <= "000000";
            when "0010110101001" => rgb <= "000000";
            when "0010110101010" => rgb <= "000000";
            when "0010110101011" => rgb <= "000000";
            when "0010110101100" => rgb <= "000000";
            when "0010110101101" => rgb <= "000000";
            when "0010110101110" => rgb <= "000000";
            when "0010110110101" => rgb <= "000000";
            when "0010110110110" => rgb <= "000000";
            when "0010110110111" => rgb <= "000000";
            when "0010110111000" => rgb <= "000000";
            when "0010110111101" => rgb <= "000000";
            when "0010110111110" => rgb <= "000000";
            when "0010110111111" => rgb <= "000000";
            when "0010111000000" => rgb <= "000000";
            when "0010111000001" => rgb <= "000000";
            when "0010111000010" => rgb <= "000000";
            when "0010111000011" => rgb <= "000000";
            when "0010111000100" => rgb <= "000000";
            when "0010111000101" => rgb <= "000000";
            when "0010111000110" => rgb <= "000000";
            when "0010111001010" => rgb <= "000000";
            when "0010111001011" => rgb <= "000000";
            when "0010111001100" => rgb <= "000000";
            when "0010111001101" => rgb <= "000000";
            when "0010111001110" => rgb <= "000000";
            when "0011000000001" => rgb <= "000000";
            when "0011000000010" => rgb <= "000000";
            when "0011000000111" => rgb <= "000000";
            when "0011000001000" => rgb <= "000000";
            when "0011000001011" => rgb <= "000000";
            when "0011000001100" => rgb <= "000000";
            when "0011000010001" => rgb <= "000000";
            when "0011000010010" => rgb <= "000000";
            when "0011000010101" => rgb <= "000000";
            when "0011000010110" => rgb <= "000000";
            when "0011000010111" => rgb <= "000000";
            when "0011000011000" => rgb <= "000000";
            when "0011000011011" => rgb <= "000000";
            when "0011000011100" => rgb <= "000000";
            when "0011000011111" => rgb <= "000000";
            when "0011000100000" => rgb <= "000000";
            when "0011000101001" => rgb <= "000000";
            when "0011000101010" => rgb <= "000000";
            when "0011000101111" => rgb <= "000000";
            when "0011000110000" => rgb <= "000000";
            when "0011000110011" => rgb <= "000000";
            when "0011000110100" => rgb <= "000000";
            when "0011000111001" => rgb <= "000000";
            when "0011000111010" => rgb <= "000000";
            when "0011001000001" => rgb <= "000000";
            when "0011001000010" => rgb <= "000000";
            when "0011001001000" => rgb <= "000000";
            when "0011001001001" => rgb <= "000000";
            when "0011010000001" => rgb <= "000000";
            when "0011010000010" => rgb <= "000000";
            when "0011010000111" => rgb <= "000000";
            when "0011010001000" => rgb <= "000000";
            when "0011010001011" => rgb <= "000000";
            when "0011010001100" => rgb <= "000000";
            when "0011010010001" => rgb <= "000000";
            when "0011010010010" => rgb <= "000000";
            when "0011010010101" => rgb <= "000000";
            when "0011010010110" => rgb <= "000000";
            when "0011010010111" => rgb <= "000000";
            when "0011010011000" => rgb <= "000000";
            when "0011010011011" => rgb <= "000000";
            when "0011010011100" => rgb <= "000000";
            when "0011010011111" => rgb <= "000000";
            when "0011010100000" => rgb <= "000000";
            when "0011010101001" => rgb <= "000000";
            when "0011010101010" => rgb <= "000000";
            when "0011010101111" => rgb <= "000000";
            when "0011010110000" => rgb <= "000000";
            when "0011010110011" => rgb <= "000000";
            when "0011010110100" => rgb <= "000000";
            when "0011010111001" => rgb <= "000000";
            when "0011010111010" => rgb <= "000000";
            when "0011011000001" => rgb <= "000000";
            when "0011011000010" => rgb <= "000000";
            when "0011011001000" => rgb <= "000000";
            when "0011011001001" => rgb <= "000000";
            when "0011100000001" => rgb <= "000000";
            when "0011100000010" => rgb <= "000000";
            when "0011100001011" => rgb <= "000000";
            when "0011100001100" => rgb <= "000000";
            when "0011100010001" => rgb <= "000000";
            when "0011100010010" => rgb <= "000000";
            when "0011100010101" => rgb <= "000000";
            when "0011100010110" => rgb <= "000000";
            when "0011100011001" => rgb <= "000000";
            when "0011100011010" => rgb <= "000000";
            when "0011100011011" => rgb <= "000000";
            when "0011100011100" => rgb <= "000000";
            when "0011100011111" => rgb <= "000000";
            when "0011100100000" => rgb <= "000000";
            when "0011100100011" => rgb <= "000000";
            when "0011100100100" => rgb <= "000000";
            when "0011100100101" => rgb <= "000000";
            when "0011100100110" => rgb <= "000000";
            when "0011100101001" => rgb <= "000000";
            when "0011100101010" => rgb <= "000000";
            when "0011100101011" => rgb <= "000000";
            when "0011100101100" => rgb <= "000000";
            when "0011100101101" => rgb <= "000000";
            when "0011100101110" => rgb <= "000000";
            when "0011100110011" => rgb <= "000000";
            when "0011100110100" => rgb <= "000000";
            when "0011100110101" => rgb <= "000000";
            when "0011100110110" => rgb <= "000000";
            when "0011100110111" => rgb <= "000000";
            when "0011100111000" => rgb <= "000000";
            when "0011100111001" => rgb <= "000000";
            when "0011100111010" => rgb <= "000000";
            when "0011101000001" => rgb <= "000000";
            when "0011101000010" => rgb <= "000000";
            when "0011101001010" => rgb <= "000000";
            when "0011101001011" => rgb <= "000000";
            when "0011101001100" => rgb <= "000000";
            when "0011101001101" => rgb <= "000000";
            when "0011110000001" => rgb <= "000000";
            when "0011110000010" => rgb <= "000000";
            when "0011110001011" => rgb <= "000000";
            when "0011110001100" => rgb <= "000000";
            when "0011110010001" => rgb <= "000000";
            when "0011110010010" => rgb <= "000000";
            when "0011110010101" => rgb <= "000000";
            when "0011110010110" => rgb <= "000000";
            when "0011110011001" => rgb <= "000000";
            when "0011110011010" => rgb <= "000000";
            when "0011110011011" => rgb <= "000000";
            when "0011110011100" => rgb <= "000000";
            when "0011110011111" => rgb <= "000000";
            when "0011110100000" => rgb <= "000000";
            when "0011110100011" => rgb <= "000000";
            when "0011110100100" => rgb <= "000000";
            when "0011110100101" => rgb <= "000000";
            when "0011110100110" => rgb <= "000000";
            when "0011110101001" => rgb <= "000000";
            when "0011110101010" => rgb <= "000000";
            when "0011110101011" => rgb <= "000000";
            when "0011110101100" => rgb <= "000000";
            when "0011110101101" => rgb <= "000000";
            when "0011110101110" => rgb <= "000000";
            when "0011110110011" => rgb <= "000000";
            when "0011110110100" => rgb <= "000000";
            when "0011110110101" => rgb <= "000000";
            when "0011110110110" => rgb <= "000000";
            when "0011110110111" => rgb <= "000000";
            when "0011110111000" => rgb <= "000000";
            when "0011110111001" => rgb <= "000000";
            when "0011110111010" => rgb <= "000000";
            when "0011111000001" => rgb <= "000000";
            when "0011111000010" => rgb <= "000000";
            when "0011111001010" => rgb <= "000000";
            when "0011111001011" => rgb <= "000000";
            when "0011111001100" => rgb <= "000000";
            when "0011111001101" => rgb <= "000000";
            when "0100000000001" => rgb <= "000000";
            when "0100000000010" => rgb <= "000000";
            when "0100000000111" => rgb <= "000000";
            when "0100000001000" => rgb <= "000000";
            when "0100000001011" => rgb <= "000000";
            when "0100000001100" => rgb <= "000000";
            when "0100000010001" => rgb <= "000000";
            when "0100000010010" => rgb <= "000000";
            when "0100000010101" => rgb <= "000000";
            when "0100000010110" => rgb <= "000000";
            when "0100000011011" => rgb <= "000000";
            when "0100000011100" => rgb <= "000000";
            when "0100000011111" => rgb <= "000000";
            when "0100000100000" => rgb <= "000000";
            when "0100000100101" => rgb <= "000000";
            when "0100000100110" => rgb <= "000000";
            when "0100000101001" => rgb <= "000000";
            when "0100000101010" => rgb <= "000000";
            when "0100000101101" => rgb <= "000000";
            when "0100000101110" => rgb <= "000000";
            when "0100000110011" => rgb <= "000000";
            when "0100000110100" => rgb <= "000000";
            when "0100000111001" => rgb <= "000000";
            when "0100000111010" => rgb <= "000000";
            when "0100001000001" => rgb <= "000000";
            when "0100001000010" => rgb <= "000000";
            when "0100001001110" => rgb <= "000000";
            when "0100010000001" => rgb <= "000000";
            when "0100010000010" => rgb <= "000000";
            when "0100010000111" => rgb <= "000000";
            when "0100010001000" => rgb <= "000000";
            when "0100010001011" => rgb <= "000000";
            when "0100010001100" => rgb <= "000000";
            when "0100010010001" => rgb <= "000000";
            when "0100010010010" => rgb <= "000000";
            when "0100010010101" => rgb <= "000000";
            when "0100010010110" => rgb <= "000000";
            when "0100010011011" => rgb <= "000000";
            when "0100010011100" => rgb <= "000000";
            when "0100010011111" => rgb <= "000000";
            when "0100010100000" => rgb <= "000000";
            when "0100010100101" => rgb <= "000000";
            when "0100010100110" => rgb <= "000000";
            when "0100010101001" => rgb <= "000000";
            when "0100010101010" => rgb <= "000000";
            when "0100010101101" => rgb <= "000000";
            when "0100010101110" => rgb <= "000000";
            when "0100010110011" => rgb <= "000000";
            when "0100010110100" => rgb <= "000000";
            when "0100010111001" => rgb <= "000000";
            when "0100010111010" => rgb <= "000000";
            when "0100011000001" => rgb <= "000000";
            when "0100011000010" => rgb <= "000000";
            when "0100011001110" => rgb <= "000000";
            when "0100100000011" => rgb <= "000000";
            when "0100100000100" => rgb <= "000000";
            when "0100100000101" => rgb <= "000000";
            when "0100100000110" => rgb <= "000000";
            when "0100100001101" => rgb <= "000000";
            when "0100100001110" => rgb <= "000000";
            when "0100100001111" => rgb <= "000000";
            when "0100100010000" => rgb <= "000000";
            when "0100100010101" => rgb <= "000000";
            when "0100100010110" => rgb <= "000000";
            when "0100100011011" => rgb <= "000000";
            when "0100100011100" => rgb <= "000000";
            when "0100100100001" => rgb <= "000000";
            when "0100100100010" => rgb <= "000000";
            when "0100100100011" => rgb <= "000000";
            when "0100100100100" => rgb <= "000000";
            when "0100100101001" => rgb <= "000000";
            when "0100100101010" => rgb <= "000000";
            when "0100100101111" => rgb <= "000000";
            when "0100100110000" => rgb <= "000000";
            when "0100100110011" => rgb <= "000000";
            when "0100100110100" => rgb <= "000000";
            when "0100100111001" => rgb <= "000000";
            when "0100100111010" => rgb <= "000000";
            when "0100101000001" => rgb <= "000000";
            when "0100101000010" => rgb <= "000000";
            when "0100101001000" => rgb <= "000000";
            when "0100101001001" => rgb <= "000000";
            when "0100101001010" => rgb <= "000000";
            when "0100101001011" => rgb <= "000000";
            when "0100101001100" => rgb <= "000000";
            when "0100101001101" => rgb <= "000000";
            when "0100110000011" => rgb <= "000000";
            when "0100110000100" => rgb <= "000000";
            when "0100110000101" => rgb <= "000000";
            when "0100110000110" => rgb <= "000000";
            when "0100110001101" => rgb <= "000000";
            when "0100110001110" => rgb <= "000000";
            when "0100110001111" => rgb <= "000000";
            when "0100110010000" => rgb <= "000000";
            when "0100110010101" => rgb <= "000000";
            when "0100110010110" => rgb <= "000000";
            when "0100110011011" => rgb <= "000000";
            when "0100110011100" => rgb <= "000000";
            when "0100110100001" => rgb <= "000000";
            when "0100110100010" => rgb <= "000000";
            when "0100110100011" => rgb <= "000000";
            when "0100110100100" => rgb <= "000000";
            when "0100110101001" => rgb <= "000000";
            when "0100110101010" => rgb <= "000000";
            when "0100110101111" => rgb <= "000000";
            when "0100110110000" => rgb <= "000000";
            when "0100110110011" => rgb <= "000000";
            when "0100110110100" => rgb <= "000000";
            when "0100110111001" => rgb <= "000000";
            when "0100110111010" => rgb <= "000000";
            when "0100111000001" => rgb <= "000000";
            when "0100111000010" => rgb <= "000000";
            when "0100111001000" => rgb <= "000000";
            when "0100111001001" => rgb <= "000000";
            when "0100111001010" => rgb <= "000000";
            when "0100111001011" => rgb <= "000000";
            when "0100111001100" => rgb <= "000000";
            when "0100111001101" => rgb <= "000000";
            when "0101110000101" => rgb <= "000000";
            when "0101110001001" => rgb <= "000000";
            when "0101110001100" => rgb <= "000000";
            when "0101110001101" => rgb <= "000000";
            when "0101110010000" => rgb <= "000000";
            when "0101110010011" => rgb <= "000000";
            when "0101110011000" => rgb <= "000000";
            when "0101110011001" => rgb <= "000000";
            when "0101110011100" => rgb <= "000000";
            when "0101110011101" => rgb <= "000000";
            when "0101110011110" => rgb <= "000000";
            when "0101110100001" => rgb <= "000000";
            when "0101110100010" => rgb <= "000000";
            when "0101110100011" => rgb <= "000000";
            when "0101110100100" => rgb <= "000000";
            when "0101110101001" => rgb <= "000000";
            when "0101110101010" => rgb <= "000000";
            when "0101110110000" => rgb <= "000000";
            when "0101110110001" => rgb <= "000000";
            when "0101110110100" => rgb <= "000000";
            when "0101110110111" => rgb <= "000000";
            when "0101110111001" => rgb <= "000000";
            when "0101110111010" => rgb <= "000000";
            when "0101110111011" => rgb <= "000000";
            when "0101110111101" => rgb <= "000000";
            when "0101110111110" => rgb <= "000000";
            when "0101110111111" => rgb <= "000000";
            when "0101111000000" => rgb <= "000000";
            when "0101111000001" => rgb <= "000000";
            when "0101111000100" => rgb <= "000000";
            when "0101111000101" => rgb <= "000000";
            when "0101111001000" => rgb <= "000000";
            when "0101111001001" => rgb <= "000000";
            when "0101111001010" => rgb <= "000000";
            when "0110000000101" => rgb <= "000000";
            when "0110000001001" => rgb <= "000000";
            when "0110000001011" => rgb <= "000000";
            when "0110000001110" => rgb <= "000000";
            when "0110000010000" => rgb <= "000000";
            when "0110000010011" => rgb <= "000000";
            when "0110000010111" => rgb <= "000000";
            when "0110000011010" => rgb <= "000000";
            when "0110000011100" => rgb <= "000000";
            when "0110000011111" => rgb <= "000000";
            when "0110000100001" => rgb <= "000000";
            when "0110000101000" => rgb <= "000000";
            when "0110000101011" => rgb <= "000000";
            when "0110000101111" => rgb <= "000000";
            when "0110000110100" => rgb <= "000000";
            when "0110000110111" => rgb <= "000000";
            when "0110000111010" => rgb <= "000000";
            when "0110000111111" => rgb <= "000000";
            when "0110001000011" => rgb <= "000000";
            when "0110001000110" => rgb <= "000000";
            when "0110001001000" => rgb <= "000000";
            when "0110001001011" => rgb <= "000000";
            when "0110010000110" => rgb <= "000000";
            when "0110010000111" => rgb <= "000000";
            when "0110010001000" => rgb <= "000000";
            when "0110010001011" => rgb <= "000000";
            when "0110010001110" => rgb <= "000000";
            when "0110010010000" => rgb <= "000000";
            when "0110010010011" => rgb <= "000000";
            when "0110010010111" => rgb <= "000000";
            when "0110010011000" => rgb <= "000000";
            when "0110010011001" => rgb <= "000000";
            when "0110010011010" => rgb <= "000000";
            when "0110010011100" => rgb <= "000000";
            when "0110010011101" => rgb <= "000000";
            when "0110010011110" => rgb <= "000000";
            when "0110010100001" => rgb <= "000000";
            when "0110010100010" => rgb <= "000000";
            when "0110010100011" => rgb <= "000000";
            when "0110010101000" => rgb <= "000000";
            when "0110010101001" => rgb <= "000000";
            when "0110010101010" => rgb <= "000000";
            when "0110010101011" => rgb <= "000000";
            when "0110010101111" => rgb <= "000000";
            when "0110010110001" => rgb <= "000000";
            when "0110010110010" => rgb <= "000000";
            when "0110010110100" => rgb <= "000000";
            when "0110010110111" => rgb <= "000000";
            when "0110010111010" => rgb <= "000000";
            when "0110010111111" => rgb <= "000000";
            when "0110011000011" => rgb <= "000000";
            when "0110011000100" => rgb <= "000000";
            when "0110011000101" => rgb <= "000000";
            when "0110011000110" => rgb <= "000000";
            when "0110011001000" => rgb <= "000000";
            when "0110011001001" => rgb <= "000000";
            when "0110011001010" => rgb <= "000000";
            when "0110100000111" => rgb <= "000000";
            when "0110100001011" => rgb <= "000000";
            when "0110100001110" => rgb <= "000000";
            when "0110100010000" => rgb <= "000000";
            when "0110100010011" => rgb <= "000000";
            when "0110100010111" => rgb <= "000000";
            when "0110100011010" => rgb <= "000000";
            when "0110100011100" => rgb <= "000000";
            when "0110100011110" => rgb <= "000000";
            when "0110100100001" => rgb <= "000000";
            when "0110100101000" => rgb <= "000000";
            when "0110100101011" => rgb <= "000000";
            when "0110100101111" => rgb <= "000000";
            when "0110100110010" => rgb <= "000000";
            when "0110100110100" => rgb <= "000000";
            when "0110100110111" => rgb <= "000000";
            when "0110100111010" => rgb <= "000000";
            when "0110100111111" => rgb <= "000000";
            when "0110101000011" => rgb <= "000000";
            when "0110101000110" => rgb <= "000000";
            when "0110101001000" => rgb <= "000000";
            when "0110101001010" => rgb <= "000000";
            when "0110110000111" => rgb <= "000000";
            when "0110110001100" => rgb <= "000000";
            when "0110110001101" => rgb <= "000000";
            when "0110110010001" => rgb <= "000000";
            when "0110110010010" => rgb <= "000000";
            when "0110110010111" => rgb <= "000000";
            when "0110110011010" => rgb <= "000000";
            when "0110110011100" => rgb <= "000000";
            when "0110110011111" => rgb <= "000000";
            when "0110110100001" => rgb <= "000000";
            when "0110110100010" => rgb <= "000000";
            when "0110110100011" => rgb <= "000000";
            when "0110110100100" => rgb <= "000000";
            when "0110110101000" => rgb <= "000000";
            when "0110110101011" => rgb <= "000000";
            when "0110110110000" => rgb <= "000000";
            when "0110110110001" => rgb <= "000000";
            when "0110110110101" => rgb <= "000000";
            when "0110110110110" => rgb <= "000000";
            when "0110110111001" => rgb <= "000000";
            when "0110110111010" => rgb <= "000000";
            when "0110110111011" => rgb <= "000000";
            when "0110110111111" => rgb <= "000000";
            when "0110111000011" => rgb <= "000000";
            when "0110111000110" => rgb <= "000000";
            when "0110111001000" => rgb <= "000000";
            when "0110111001011" => rgb <= "000000";
            when "0111100011010" => rgb <= "000000";
            when "0111100011101" => rgb <= "000000";
            when "0111100011111" => rgb <= "000000";
            when "0111100100000" => rgb <= "000000";
            when "0111100100001" => rgb <= "000000";
            when "0111100100010" => rgb <= "000000";
            when "0111100100100" => rgb <= "000000";
            when "0111100100101" => rgb <= "000000";
            when "0111100100110" => rgb <= "000000";
            when "0111100101010" => rgb <= "000000";
            when "0111100101011" => rgb <= "000000";
            when "0111100101111" => rgb <= "000000";
            when "0111100110011" => rgb <= "000000";
            when "0111110011010" => rgb <= "000000";
            when "0111110011101" => rgb <= "000000";
            when "0111110011111" => rgb <= "000000";
            when "0111110100100" => rgb <= "000000";
            when "0111110100111" => rgb <= "000000";
            when "0111110101001" => rgb <= "000000";
            when "0111110101100" => rgb <= "000000";
            when "0111110101111" => rgb <= "000000";
            when "0111110110011" => rgb <= "000000";
            when "1000000011010" => rgb <= "000000";
            when "1000000011011" => rgb <= "000000";
            when "1000000011100" => rgb <= "000000";
            when "1000000011101" => rgb <= "000000";
            when "1000000011111" => rgb <= "000000";
            when "1000000100000" => rgb <= "000000";
            when "1000000100001" => rgb <= "000000";
            when "1000000100100" => rgb <= "000000";
            when "1000000100101" => rgb <= "000000";
            when "1000000100110" => rgb <= "000000";
            when "1000000101001" => rgb <= "000000";
            when "1000000101100" => rgb <= "000000";
            when "1000000101111" => rgb <= "000000";
            when "1000000110011" => rgb <= "000000";
            when "1000010011010" => rgb <= "000000";
            when "1000010011101" => rgb <= "000000";
            when "1000010011111" => rgb <= "000000";
            when "1000010100100" => rgb <= "000000";
            when "1000010100110" => rgb <= "000000";
            when "1000010101001" => rgb <= "000000";
            when "1000010101100" => rgb <= "000000";
            when "1000100011010" => rgb <= "000000";
            when "1000100011101" => rgb <= "000000";
            when "1000100011111" => rgb <= "000000";
            when "1000100100000" => rgb <= "000000";
            when "1000100100001" => rgb <= "000000";
            when "1000100100010" => rgb <= "000000";
            when "1000100100100" => rgb <= "000000";
            when "1000100100111" => rgb <= "000000";
            when "1000100101010" => rgb <= "000000";
            when "1000100101011" => rgb <= "000000";
            when "1000100101111" => rgb <= "000000";
            when "1000100110011" => rgb <= "000000";
            when "1001010001110" => rgb <= "000000";
            when "1001010001111" => rgb <= "000000";
            when "1001010010000" => rgb <= "000000";
            when "1001010010011" => rgb <= "000000";
            when "1001010010100" => rgb <= "000000";
            when "1001010011000" => rgb <= "000000";
            when "1001010011001" => rgb <= "000000";
            when "1001010011100" => rgb <= "000000";
            when "1001010011101" => rgb <= "000000";
            when "1001010011110" => rgb <= "000000";
            when "1001010100001" => rgb <= "000000";
            when "1001010100010" => rgb <= "000000";
            when "1001010100011" => rgb <= "000000";
            when "1001010100100" => rgb <= "000000";
            when "1001100001101" => rgb <= "000000";
            when "1001100010010" => rgb <= "000000";
            when "1001100010101" => rgb <= "000000";
            when "1001100010111" => rgb <= "000000";
            when "1001100011010" => rgb <= "000000";
            when "1001100011100" => rgb <= "000000";
            when "1001100011111" => rgb <= "000000";
            when "1001100100001" => rgb <= "000000";
            when "1001100100111" => rgb <= "000000";
            when "1001110001110" => rgb <= "000000";
            when "1001110001111" => rgb <= "000000";
            when "1001110010010" => rgb <= "000000";
            when "1001110010111" => rgb <= "000000";
            when "1001110011010" => rgb <= "000000";
            when "1001110011100" => rgb <= "000000";
            when "1001110011101" => rgb <= "000000";
            when "1001110011110" => rgb <= "000000";
            when "1001110100001" => rgb <= "000000";
            when "1001110100010" => rgb <= "000000";
            when "1001110100011" => rgb <= "000000";
            when "1010000010000" => rgb <= "000000";
            when "1010000010010" => rgb <= "000000";
            when "1010000010101" => rgb <= "000000";
            when "1010000010111" => rgb <= "000000";
            when "1010000011010" => rgb <= "000000";
            when "1010000011100" => rgb <= "000000";
            when "1010000011110" => rgb <= "000000";
            when "1010000100001" => rgb <= "000000";
            when "1010000100111" => rgb <= "000000";
            when "1010010001101" => rgb <= "000000";
            when "1010010001110" => rgb <= "000000";
            when "1010010001111" => rgb <= "000000";
            when "1010010010011" => rgb <= "000000";
            when "1010010010100" => rgb <= "000000";
            when "1010010011000" => rgb <= "000000";
            when "1010010011001" => rgb <= "000000";
            when "1010010011100" => rgb <= "000000";
            when "1010010011111" => rgb <= "000000";
            when "1010010100001" => rgb <= "000000";
            when "1010010100010" => rgb <= "000000";
            when "1010010100011" => rgb <= "000000";
            when "1010010100100" => rgb <= "000000";
            when "1010010111011" => rgb <= "100000";
            when "1010010111100" => rgb <= "100000";
            when "1010010111101" => rgb <= "100000";
            when "1010010111110" => rgb <= "100000";
            when "1010010111111" => rgb <= "100000";
            when "1010011000000" => rgb <= "100000";
            when "1010011000001" => rgb <= "100000";
            when "1010011000010" => rgb <= "100000";
            when "1010011000011" => rgb <= "100000";
            when "1010011000100" => rgb <= "100000";
            when "1010011000110" => rgb <= "100000";
            when "1010011000111" => rgb <= "100000";
            when "1010011001000" => rgb <= "100000";
            when "1010100111001" => rgb <= "100000";
            when "1010100111010" => rgb <= "100000";
            when "1010100111011" => rgb <= "100000";
            when "1010100111100" => rgb <= "100000";
            when "1010100111101" => rgb <= "100000";
            when "1010100111110" => rgb <= "100000";
            when "1010100111111" => rgb <= "100000";
            when "1010101000000" => rgb <= "100000";
            when "1010101000001" => rgb <= "100000";
            when "1010101000010" => rgb <= "100000";
            when "1010101000011" => rgb <= "110100";
            when "1010101000100" => rgb <= "100000";
            when "1010101000101" => rgb <= "100000";
            when "1010101000110" => rgb <= "100000";
            when "1010101000111" => rgb <= "110100";
            when "1010101001000" => rgb <= "100000";
            when "1010101001001" => rgb <= "100000";
            when "1010101001010" => rgb <= "100000";
            when "1010110001001" => rgb <= "010000";
            when "1010110001010" => rgb <= "010000";
            when "1010110001011" => rgb <= "010000";
            when "1010110001100" => rgb <= "010000";
            when "1010110001101" => rgb <= "010000";
            when "1010110001110" => rgb <= "010000";
            when "1010110001111" => rgb <= "010000";
            when "1010110011010" => rgb <= "010000";
            when "1010110011011" => rgb <= "010000";
            when "1010110011100" => rgb <= "010000";
            when "1010110011101" => rgb <= "010000";
            when "1010110011110" => rgb <= "010000";
            when "1010110011111" => rgb <= "010000";
            when "1010110100000" => rgb <= "010000";
            when "1010110110101" => rgb <= "100000";
            when "1010110110110" => rgb <= "100000";
            when "1010110110111" => rgb <= "100000";
            when "1010110111000" => rgb <= "100000";
            when "1010110111001" => rgb <= "100000";
            when "1010110111010" => rgb <= "100000";
            when "1010110111011" => rgb <= "100000";
            when "1010110111100" => rgb <= "100000";
            when "1010110111101" => rgb <= "110100";
            when "1010110111110" => rgb <= "110100";
            when "1010110111111" => rgb <= "110100";
            when "1010111000000" => rgb <= "100000";
            when "1010111000001" => rgb <= "100000";
            when "1010111000010" => rgb <= "110100";
            when "1010111000011" => rgb <= "110100";
            when "1010111000100" => rgb <= "100000";
            when "1010111000101" => rgb <= "110100";
            when "1010111000110" => rgb <= "110100";
            when "1010111000111" => rgb <= "110100";
            when "1010111001000" => rgb <= "110100";
            when "1010111001001" => rgb <= "110100";
            when "1010111001010" => rgb <= "100000";
            when "1010111001011" => rgb <= "100000";
            when "1010111001100" => rgb <= "100000";
            when "1011000001000" => rgb <= "010000";
            when "1011000001001" => rgb <= "010000";
            when "1011000001010" => rgb <= "010000";
            when "1011000001011" => rgb <= "010000";
            when "1011000001100" => rgb <= "010000";
            when "1011000001101" => rgb <= "010000";
            when "1011000001110" => rgb <= "010000";
            when "1011000001111" => rgb <= "010000";
            when "1011000010000" => rgb <= "010000";
            when "1011000010001" => rgb <= "010000";
            when "1011000010010" => rgb <= "010000";
            when "1011000010011" => rgb <= "010000";
            when "1011000010100" => rgb <= "010000";
            when "1011000011000" => rgb <= "010000";
            when "1011000011001" => rgb <= "010000";
            when "1011000011010" => rgb <= "010000";
            when "1011000011011" => rgb <= "010000";
            when "1011000011100" => rgb <= "010000";
            when "1011000011101" => rgb <= "010000";
            when "1011000011110" => rgb <= "010000";
            when "1011000011111" => rgb <= "010000";
            when "1011000100000" => rgb <= "010000";
            when "1011000100001" => rgb <= "010000";
            when "1011000100010" => rgb <= "010000";
            when "1011000100011" => rgb <= "010000";
            when "1011000110100" => rgb <= "100000";
            when "1011000110101" => rgb <= "100000";
            when "1011000110110" => rgb <= "100000";
            when "1011000110111" => rgb <= "100000";
            when "1011000111000" => rgb <= "100000";
            when "1011000111001" => rgb <= "100000";
            when "1011000111010" => rgb <= "110100";
            when "1011000111011" => rgb <= "110100";
            when "1011000111100" => rgb <= "110100";
            when "1011000111101" => rgb <= "110100";
            when "1011000111110" => rgb <= "110100";
            when "1011000111111" => rgb <= "110100";
            when "1011001000000" => rgb <= "110100";
            when "1011001000001" => rgb <= "100000";
            when "1011001000010" => rgb <= "110100";
            when "1011001000011" => rgb <= "110100";
            when "1011001000100" => rgb <= "110100";
            when "1011001000101" => rgb <= "110100";
            when "1011001000110" => rgb <= "110100";
            when "1011001000111" => rgb <= "110100";
            when "1011001001000" => rgb <= "100000";
            when "1011001001001" => rgb <= "100000";
            when "1011001001010" => rgb <= "100000";
            when "1011010000111" => rgb <= "010000";
            when "1011010001000" => rgb <= "010000";
            when "1011010001001" => rgb <= "010000";
            when "1011010001010" => rgb <= "010000";
            when "1011010001011" => rgb <= "010000";
            when "1011010001100" => rgb <= "010000";
            when "1011010001101" => rgb <= "010000";
            when "1011010001110" => rgb <= "010000";
            when "1011010001111" => rgb <= "010000";
            when "1011010010000" => rgb <= "010000";
            when "1011010010001" => rgb <= "010000";
            when "1011010010010" => rgb <= "010000";
            when "1011010010011" => rgb <= "010000";
            when "1011010010100" => rgb <= "010000";
            when "1011010010101" => rgb <= "010000";
            when "1011010010110" => rgb <= "010000";
            when "1011010010111" => rgb <= "010000";
            when "1011010011000" => rgb <= "010000";
            when "1011010011101" => rgb <= "010000";
            when "1011010011110" => rgb <= "010000";
            when "1011010011111" => rgb <= "010000";
            when "1011010100000" => rgb <= "010000";
            when "1011010100001" => rgb <= "010000";
            when "1011010100010" => rgb <= "010000";
            when "1011010100011" => rgb <= "010000";
            when "1011010110010" => rgb <= "100000";
            when "1011010110011" => rgb <= "100000";
            when "1011010110100" => rgb <= "100000";
            when "1011010110101" => rgb <= "100000";
            when "1011010110110" => rgb <= "100000";
            when "1011010110111" => rgb <= "000000";
            when "1011010111000" => rgb <= "100000";
            when "1011010111001" => rgb <= "110100";
            when "1011010111010" => rgb <= "110100";
            when "1011010111011" => rgb <= "110100";
            when "1011010111100" => rgb <= "110100";
            when "1011010111101" => rgb <= "110100";
            when "1011010111110" => rgb <= "110100";
            when "1011010111111" => rgb <= "110100";
            when "1011011000000" => rgb <= "110100";
            when "1011011000001" => rgb <= "110100";
            when "1011011000010" => rgb <= "110100";
            when "1011011000011" => rgb <= "110100";
            when "1011011000100" => rgb <= "110100";
            when "1011011000101" => rgb <= "110100";
            when "1011011000110" => rgb <= "110100";
            when "1011011000111" => rgb <= "100000";
            when "1011011001000" => rgb <= "100000";
            when "1011011001001" => rgb <= "100000";
            when "1011100000110" => rgb <= "010000";
            when "1011100000111" => rgb <= "010000";
            when "1011100001000" => rgb <= "010000";
            when "1011100001001" => rgb <= "000000";
            when "1011100001010" => rgb <= "000000";
            when "1011100001011" => rgb <= "010000";
            when "1011100001100" => rgb <= "000000";
            when "1011100001101" => rgb <= "010000";
            when "1011100010010" => rgb <= "010000";
            when "1011100010011" => rgb <= "010000";
            when "1011100010100" => rgb <= "010000";
            when "1011100010101" => rgb <= "010000";
            when "1011100010110" => rgb <= "010000";
            when "1011100011111" => rgb <= "010000";
            when "1011100100000" => rgb <= "010000";
            when "1011100100001" => rgb <= "010000";
            when "1011100110001" => rgb <= "100000";
            when "1011100110010" => rgb <= "100000";
            when "1011100110011" => rgb <= "100000";
            when "1011100110100" => rgb <= "000000";
            when "1011100110101" => rgb <= "100000";
            when "1011100110110" => rgb <= "010000";
            when "1011100110111" => rgb <= "010000";
            when "1011100111000" => rgb <= "110100";
            when "1011100111001" => rgb <= "110100";
            when "1011100111010" => rgb <= "110100";
            when "1011100111011" => rgb <= "110100";
            when "1011100111100" => rgb <= "111000";
            when "1011100111101" => rgb <= "111000";
            when "1011100111110" => rgb <= "111000";
            when "1011100111111" => rgb <= "110100";
            when "1011101000000" => rgb <= "110100";
            when "1011101000001" => rgb <= "110100";
            when "1011101000010" => rgb <= "110100";
            when "1011101000011" => rgb <= "110100";
            when "1011101000100" => rgb <= "110100";
            when "1011101000101" => rgb <= "100000";
            when "1011101000110" => rgb <= "100000";
            when "1011101000111" => rgb <= "100000";
            when "1011101001000" => rgb <= "100000";
            when "1011101001001" => rgb <= "100000";
            when "1011110000110" => rgb <= "010000";
            when "1011110000111" => rgb <= "010000";
            when "1011110001000" => rgb <= "010000";
            when "1011110001001" => rgb <= "000000";
            when "1011110001010" => rgb <= "000000";
            when "1011110001011" => rgb <= "010000";
            when "1011110001100" => rgb <= "010000";
            when "1011110001101" => rgb <= "010000";
            when "1011110001110" => rgb <= "010000";
            when "1011110011101" => rgb <= "010000";
            when "1011110011110" => rgb <= "010000";
            when "1011110011111" => rgb <= "010000";
            when "1011110100000" => rgb <= "010000";
            when "1011110101111" => rgb <= "100000";
            when "1011110110000" => rgb <= "100000";
            when "1011110110001" => rgb <= "100000";
            when "1011110110010" => rgb <= "100000";
            when "1011110110011" => rgb <= "010000";
            when "1011110110100" => rgb <= "010000";
            when "1011110110101" => rgb <= "010000";
            when "1011110110110" => rgb <= "010000";
            when "1011110110111" => rgb <= "010000";
            when "1011110111000" => rgb <= "110100";
            when "1011110111001" => rgb <= "110100";
            when "1011110111010" => rgb <= "110100";
            when "1011110111011" => rgb <= "110100";
            when "1011110111100" => rgb <= "111000";
            when "1011110111101" => rgb <= "111000";
            when "1011110111110" => rgb <= "111000";
            when "1011110111111" => rgb <= "111000";
            when "1011111000000" => rgb <= "111000";
            when "1011111000001" => rgb <= "110100";
            when "1011111000010" => rgb <= "110100";
            when "1011111000011" => rgb <= "110100";
            when "1011111000100" => rgb <= "110100";
            when "1011111000101" => rgb <= "110100";
            when "1011111000110" => rgb <= "100000";
            when "1011111000111" => rgb <= "100000";
            when "1011111001000" => rgb <= "100000";
            when "1100000000110" => rgb <= "010000";
            when "1100000000111" => rgb <= "010000";
            when "1100000001000" => rgb <= "010000";
            when "1100000001001" => rgb <= "000000";
            when "1100000001010" => rgb <= "000000";
            when "1100000001011" => rgb <= "010000";
            when "1100000001100" => rgb <= "000000";
            when "1100000001101" => rgb <= "010000";
            when "1100000001110" => rgb <= "010000";
            when "1100000011100" => rgb <= "010000";
            when "1100000011101" => rgb <= "010000";
            when "1100000011110" => rgb <= "010000";
            when "1100000101111" => rgb <= "100000";
            when "1100000110000" => rgb <= "100000";
            when "1100000110001" => rgb <= "100000";
            when "1100000110010" => rgb <= "010000";
            when "1100000110011" => rgb <= "010000";
            when "1100000110100" => rgb <= "000000";
            when "1100000110101" => rgb <= "010000";
            when "1100000110110" => rgb <= "010000";
            when "1100000110111" => rgb <= "000000";
            when "1100000111000" => rgb <= "010000";
            when "1100000111001" => rgb <= "110100";
            when "1100000111010" => rgb <= "000000";
            when "1100000111011" => rgb <= "000000";
            when "1100000111100" => rgb <= "111000";
            when "1100000111101" => rgb <= "111000";
            when "1100000111110" => rgb <= "111000";
            when "1100000111111" => rgb <= "111000";
            when "1100001000000" => rgb <= "111000";
            when "1100001000001" => rgb <= "111000";
            when "1100001000010" => rgb <= "111000";
            when "1100001000011" => rgb <= "111000";
            when "1100001000100" => rgb <= "110100";
            when "1100001000101" => rgb <= "110100";
            when "1100001000110" => rgb <= "110100";
            when "1100001000111" => rgb <= "110100";
            when "1100001001000" => rgb <= "100000";
            when "1100001001001" => rgb <= "100000";
            when "1100001001010" => rgb <= "100000";
            when "1100010000110" => rgb <= "010000";
            when "1100010000111" => rgb <= "010000";
            when "1100010001000" => rgb <= "010000";
            when "1100010001001" => rgb <= "000000";
            when "1100010001010" => rgb <= "000000";
            when "1100010001011" => rgb <= "010000";
            when "1100010001100" => rgb <= "010000";
            when "1100010001101" => rgb <= "010000";
            when "1100010010110" => rgb <= "000000";
            when "1100010011100" => rgb <= "010000";
            when "1100010011101" => rgb <= "010000";
            when "1100010011110" => rgb <= "010100";
            when "1100010011111" => rgb <= "010100";
            when "1100010100000" => rgb <= "010100";
            when "1100010100001" => rgb <= "010100";
            when "1100010100010" => rgb <= "010100";
            when "1100010100011" => rgb <= "010100";
            when "1100010100100" => rgb <= "010100";
            when "1100010100101" => rgb <= "010100";
            when "1100010100110" => rgb <= "010100";
            when "1100010100111" => rgb <= "010100";
            when "1100010101000" => rgb <= "000000";
            when "1100010101001" => rgb <= "010100";
            when "1100010101010" => rgb <= "010100";
            when "1100010101011" => rgb <= "010100";
            when "1100010101100" => rgb <= "010100";
            when "1100010101101" => rgb <= "010100";
            when "1100010101110" => rgb <= "010100";
            when "1100010101111" => rgb <= "010100";
            when "1100010110000" => rgb <= "010100";
            when "1100010110001" => rgb <= "010100";
            when "1100010110010" => rgb <= "010000";
            when "1100010110011" => rgb <= "010000";
            when "1100010110100" => rgb <= "010000";
            when "1100010110101" => rgb <= "010000";
            when "1100010110110" => rgb <= "010000";
            when "1100010110111" => rgb <= "010000";
            when "1100010111000" => rgb <= "010000";
            when "1100010111001" => rgb <= "010000";
            when "1100010111010" => rgb <= "010000";
            when "1100010111011" => rgb <= "010000";
            when "1100010111100" => rgb <= "111000";
            when "1100010111101" => rgb <= "111000";
            when "1100010111110" => rgb <= "111000";
            when "1100010111111" => rgb <= "111000";
            when "1100011000000" => rgb <= "111000";
            when "1100011000001" => rgb <= "111000";
            when "1100011000010" => rgb <= "111000";
            when "1100011000011" => rgb <= "111000";
            when "1100011000100" => rgb <= "110100";
            when "1100011000101" => rgb <= "110100";
            when "1100011000110" => rgb <= "110100";
            when "1100011000111" => rgb <= "110100";
            when "1100011001000" => rgb <= "110100";
            when "1100011001001" => rgb <= "110100";
            when "1100011001010" => rgb <= "100000";
            when "1100011001011" => rgb <= "100000";
            when "1100100000110" => rgb <= "010000";
            when "1100100000111" => rgb <= "010000";
            when "1100100001000" => rgb <= "010000";
            when "1100100001001" => rgb <= "000000";
            when "1100100001010" => rgb <= "000000";
            when "1100100001011" => rgb <= "010000";
            when "1100100001100" => rgb <= "000000";
            when "1100100001101" => rgb <= "010000";
            when "1100100001110" => rgb <= "010000";
            when "1100100011100" => rgb <= "010000";
            when "1100100011101" => rgb <= "010100";
            when "1100100011110" => rgb <= "010100";
            when "1100100011111" => rgb <= "000000";
            when "1100100100000" => rgb <= "010100";
            when "1100100100001" => rgb <= "010100";
            when "1100100100010" => rgb <= "010100";
            when "1100100100011" => rgb <= "000000";
            when "1100100100100" => rgb <= "010100";
            when "1100100100101" => rgb <= "010100";
            when "1100100100110" => rgb <= "000000";
            when "1100100100111" => rgb <= "010100";
            when "1100100101000" => rgb <= "010100";
            when "1100100101001" => rgb <= "010100";
            when "1100100101010" => rgb <= "000000";
            when "1100100101011" => rgb <= "010100";
            when "1100100101100" => rgb <= "010100";
            when "1100100101101" => rgb <= "010100";
            when "1100100101110" => rgb <= "000000";
            when "1100100101111" => rgb <= "010100";
            when "1100100110000" => rgb <= "010100";
            when "1100100110001" => rgb <= "010100";
            when "1100100110010" => rgb <= "010000";
            when "1100100110011" => rgb <= "010000";
            when "1100100110100" => rgb <= "010000";
            when "1100100110101" => rgb <= "010000";
            when "1100100110110" => rgb <= "010000";
            when "1100100110111" => rgb <= "010000";
            when "1100100111000" => rgb <= "010000";
            when "1100100111001" => rgb <= "010000";
            when "1100100111010" => rgb <= "000000";
            when "1100100111011" => rgb <= "010000";
            when "1100100111100" => rgb <= "010000";
            when "1100100111101" => rgb <= "010000";
            when "1100100111110" => rgb <= "111000";
            when "1100100111111" => rgb <= "111000";
            when "1100101000000" => rgb <= "111000";
            when "1100101000001" => rgb <= "111000";
            when "1100101000010" => rgb <= "111000";
            when "1100101000011" => rgb <= "111000";
            when "1100101000100" => rgb <= "110100";
            when "1100101000101" => rgb <= "110100";
            when "1100101000110" => rgb <= "110100";
            when "1100101000111" => rgb <= "110100";
            when "1100101001000" => rgb <= "110100";
            when "1100101001001" => rgb <= "110100";
            when "1100101001010" => rgb <= "110100";
            when "1100101001011" => rgb <= "100000";
            when "1100101001100" => rgb <= "100000";
            when "1100110000110" => rgb <= "010000";
            when "1100110000111" => rgb <= "010000";
            when "1100110001000" => rgb <= "010000";
            when "1100110001001" => rgb <= "010000";
            when "1100110001010" => rgb <= "010000";
            when "1100110001011" => rgb <= "010000";
            when "1100110001100" => rgb <= "010000";
            when "1100110001101" => rgb <= "000000";
            when "1100110001110" => rgb <= "010000";
            when "1100110010110" => rgb <= "000000";
            when "1100110011100" => rgb <= "010000";
            when "1100110011101" => rgb <= "010100";
            when "1100110011110" => rgb <= "010100";
            when "1100110011111" => rgb <= "000000";
            when "1100110100000" => rgb <= "010100";
            when "1100110100001" => rgb <= "010100";
            when "1100110100010" => rgb <= "010100";
            when "1100110100011" => rgb <= "000000";
            when "1100110100100" => rgb <= "010100";
            when "1100110100101" => rgb <= "010100";
            when "1100110100110" => rgb <= "000000";
            when "1100110100111" => rgb <= "010100";
            when "1100110101000" => rgb <= "010100";
            when "1100110101001" => rgb <= "010100";
            when "1100110101010" => rgb <= "000000";
            when "1100110101011" => rgb <= "010100";
            when "1100110101100" => rgb <= "010100";
            when "1100110101101" => rgb <= "010100";
            when "1100110101110" => rgb <= "000000";
            when "1100110101111" => rgb <= "010100";
            when "1100110110000" => rgb <= "010100";
            when "1100110110001" => rgb <= "010100";
            when "1100110110010" => rgb <= "010000";
            when "1100110110011" => rgb <= "010000";
            when "1100110110100" => rgb <= "000000";
            when "1100110110101" => rgb <= "010000";
            when "1100110110110" => rgb <= "010000";
            when "1100110110111" => rgb <= "000000";
            when "1100110111000" => rgb <= "010000";
            when "1100110111001" => rgb <= "010000";
            when "1100110111010" => rgb <= "010000";
            when "1100110111011" => rgb <= "010000";
            when "1100110111100" => rgb <= "010000";
            when "1100110111101" => rgb <= "010000";
            when "1100110111110" => rgb <= "111000";
            when "1100110111111" => rgb <= "111000";
            when "1100111000000" => rgb <= "111000";
            when "1100111000001" => rgb <= "111000";
            when "1100111000010" => rgb <= "111000";
            when "1100111000011" => rgb <= "110100";
            when "1100111000100" => rgb <= "110100";
            when "1100111000101" => rgb <= "110100";
            when "1100111000110" => rgb <= "110100";
            when "1100111000111" => rgb <= "100000";
            when "1100111001000" => rgb <= "100000";
            when "1100111001001" => rgb <= "100000";
            when "1100111001010" => rgb <= "100000";
            when "1100111001011" => rgb <= "100000";
            when "1100111001100" => rgb <= "100000";
            when "1100111001101" => rgb <= "100000";
            when "1101000000110" => rgb <= "010000";
            when "1101000000111" => rgb <= "010000";
            when "1101000001000" => rgb <= "010000";
            when "1101000001001" => rgb <= "010000";
            when "1101000001010" => rgb <= "010000";
            when "1101000001011" => rgb <= "010000";
            when "1101000001100" => rgb <= "010000";
            when "1101000001101" => rgb <= "000000";
            when "1101000001110" => rgb <= "010000";
            when "1101000011100" => rgb <= "010000";
            when "1101000011101" => rgb <= "010000";
            when "1101000011110" => rgb <= "010100";
            when "1101000011111" => rgb <= "010100";
            when "1101000100000" => rgb <= "010100";
            when "1101000100001" => rgb <= "010100";
            when "1101000100010" => rgb <= "010100";
            when "1101000100011" => rgb <= "010100";
            when "1101000100100" => rgb <= "010100";
            when "1101000100101" => rgb <= "010100";
            when "1101000100110" => rgb <= "010100";
            when "1101000100111" => rgb <= "010100";
            when "1101000101000" => rgb <= "000000";
            when "1101000101001" => rgb <= "010100";
            when "1101000101010" => rgb <= "010100";
            when "1101000101011" => rgb <= "010100";
            when "1101000101100" => rgb <= "010100";
            when "1101000101101" => rgb <= "010100";
            when "1101000101110" => rgb <= "010100";
            when "1101000101111" => rgb <= "010100";
            when "1101000110000" => rgb <= "010100";
            when "1101000110001" => rgb <= "010100";
            when "1101000110010" => rgb <= "010100";
            when "1101000110011" => rgb <= "010000";
            when "1101000110100" => rgb <= "010000";
            when "1101000110101" => rgb <= "010000";
            when "1101000110110" => rgb <= "010000";
            when "1101000110111" => rgb <= "010000";
            when "1101000111000" => rgb <= "010000";
            when "1101000111001" => rgb <= "010000";
            when "1101000111010" => rgb <= "010000";
            when "1101000111011" => rgb <= "010000";
            when "1101000111100" => rgb <= "010000";
            when "1101000111101" => rgb <= "010000";
            when "1101000111110" => rgb <= "111000";
            when "1101000111111" => rgb <= "111000";
            when "1101001000000" => rgb <= "111000";
            when "1101001000001" => rgb <= "110100";
            when "1101001000010" => rgb <= "110100";
            when "1101001000011" => rgb <= "110100";
            when "1101001000100" => rgb <= "110100";
            when "1101001000101" => rgb <= "100000";
            when "1101001000110" => rgb <= "100000";
            when "1101001000111" => rgb <= "100000";
            when "1101001001000" => rgb <= "100000";
            when "1101010000110" => rgb <= "010000";
            when "1101010000111" => rgb <= "010000";
            when "1101010001000" => rgb <= "010000";
            when "1101010001001" => rgb <= "010000";
            when "1101010001010" => rgb <= "010000";
            when "1101010001011" => rgb <= "000000";
            when "1101010001100" => rgb <= "010000";
            when "1101010001101" => rgb <= "000000";
            when "1101010001110" => rgb <= "010000";
            when "1101010010010" => rgb <= "010000";
            when "1101010010011" => rgb <= "010000";
            when "1101010010100" => rgb <= "010000";
            when "1101010010101" => rgb <= "010000";
            when "1101010010110" => rgb <= "010000";
            when "1101010010111" => rgb <= "010000";
            when "1101010011100" => rgb <= "010000";
            when "1101010011101" => rgb <= "010000";
            when "1101010011110" => rgb <= "010000";
            when "1101010011111" => rgb <= "010000";
            when "1101010110010" => rgb <= "100000";
            when "1101010110011" => rgb <= "100000";
            when "1101010110100" => rgb <= "000000";
            when "1101010110101" => rgb <= "100000";
            when "1101010110110" => rgb <= "100000";
            when "1101010110111" => rgb <= "010000";
            when "1101010111000" => rgb <= "010000";
            when "1101010111001" => rgb <= "010000";
            when "1101010111010" => rgb <= "000000";
            when "1101010111011" => rgb <= "010000";
            when "1101010111100" => rgb <= "010000";
            when "1101010111101" => rgb <= "010000";
            when "1101010111110" => rgb <= "111000";
            when "1101010111111" => rgb <= "111000";
            when "1101011000000" => rgb <= "110100";
            when "1101011000001" => rgb <= "110100";
            when "1101011000010" => rgb <= "110100";
            when "1101011000011" => rgb <= "100000";
            when "1101011000100" => rgb <= "100000";
            when "1101011000101" => rgb <= "100000";
            when "1101011000110" => rgb <= "100000";
            when "1101011000111" => rgb <= "100000";
            when "1101100000111" => rgb <= "010000";
            when "1101100001000" => rgb <= "010000";
            when "1101100001001" => rgb <= "010000";
            when "1101100001010" => rgb <= "010000";
            when "1101100001011" => rgb <= "000000";
            when "1101100001100" => rgb <= "010000";
            when "1101100010001" => rgb <= "010000";
            when "1101100010010" => rgb <= "010000";
            when "1101100010011" => rgb <= "010000";
            when "1101100010100" => rgb <= "010000";
            when "1101100010101" => rgb <= "010000";
            when "1101100010110" => rgb <= "010000";
            when "1101100010111" => rgb <= "010000";
            when "1101100011000" => rgb <= "010000";
            when "1101100011001" => rgb <= "010000";
            when "1101100011110" => rgb <= "010000";
            when "1101100011111" => rgb <= "010000";
            when "1101100100000" => rgb <= "010000";
            when "1101100100001" => rgb <= "010000";
            when "1101100110010" => rgb <= "100000";
            when "1101100110011" => rgb <= "100000";
            when "1101100110100" => rgb <= "100000";
            when "1101100110101" => rgb <= "100000";
            when "1101100110110" => rgb <= "100000";
            when "1101100110111" => rgb <= "000000";
            when "1101100111000" => rgb <= "010000";
            when "1101100111001" => rgb <= "010000";
            when "1101100111010" => rgb <= "010000";
            when "1101100111011" => rgb <= "010000";
            when "1101100111100" => rgb <= "110100";
            when "1101100111101" => rgb <= "110100";
            when "1101100111110" => rgb <= "110100";
            when "1101100111111" => rgb <= "110100";
            when "1101101000000" => rgb <= "110100";
            when "1101101000001" => rgb <= "110100";
            when "1101101000010" => rgb <= "110100";
            when "1101101000011" => rgb <= "100000";
            when "1101101000100" => rgb <= "100000";
            when "1101101000101" => rgb <= "100000";
            when "1101101000110" => rgb <= "100000";
            when "1101110001000" => rgb <= "010000";
            when "1101110001001" => rgb <= "010000";
            when "1101110001010" => rgb <= "010000";
            when "1101110001011" => rgb <= "010000";
            when "1101110001100" => rgb <= "010000";
            when "1101110001101" => rgb <= "010000";
            when "1101110001110" => rgb <= "010000";
            when "1101110001111" => rgb <= "010000";
            when "1101110010000" => rgb <= "010000";
            when "1101110010001" => rgb <= "010000";
            when "1101110010010" => rgb <= "010000";
            when "1101110010011" => rgb <= "010000";
            when "1101110010110" => rgb <= "010000";
            when "1101110010111" => rgb <= "010000";
            when "1101110011000" => rgb <= "010000";
            when "1101110011001" => rgb <= "010000";
            when "1101110011010" => rgb <= "010000";
            when "1101110011011" => rgb <= "010000";
            when "1101110011110" => rgb <= "010000";
            when "1101110011111" => rgb <= "010000";
            when "1101110100000" => rgb <= "010000";
            when "1101110100001" => rgb <= "010000";
            when "1101110100010" => rgb <= "010000";
            when "1101110110101" => rgb <= "100000";
            when "1101110110110" => rgb <= "100000";
            when "1101110110111" => rgb <= "100000";
            when "1101110111000" => rgb <= "100000";
            when "1101110111001" => rgb <= "100000";
            when "1101110111010" => rgb <= "000000";
            when "1101110111011" => rgb <= "000000";
            when "1101110111100" => rgb <= "100000";
            when "1101110111101" => rgb <= "100000";
            when "1101110111110" => rgb <= "100000";
            when "1101110111111" => rgb <= "110100";
            when "1101111000000" => rgb <= "110100";
            when "1101111000001" => rgb <= "100000";
            when "1101111000010" => rgb <= "100000";
            when "1101111000011" => rgb <= "100000";
            when "1101111000100" => rgb <= "100000";
            when "1101111000101" => rgb <= "100000";
            when "1101111000110" => rgb <= "100000";
            when "1110000001001" => rgb <= "010000";
            when "1110000001010" => rgb <= "010000";
            when "1110000001011" => rgb <= "010000";
            when "1110000001100" => rgb <= "010000";
            when "1110000001101" => rgb <= "010000";
            when "1110000001110" => rgb <= "010000";
            when "1110000001111" => rgb <= "010000";
            when "1110000010000" => rgb <= "010000";
            when "1110000011001" => rgb <= "010000";
            when "1110000011010" => rgb <= "010000";
            when "1110000011011" => rgb <= "010000";
            when "1110000011100" => rgb <= "010000";
            when "1110000011101" => rgb <= "010000";
            when "1110000011110" => rgb <= "010000";
            when "1110000011111" => rgb <= "010000";
            when "1110000100000" => rgb <= "010000";
            when "1110000100001" => rgb <= "010000";
            when "1110000100010" => rgb <= "010000";
            when "1110000110111" => rgb <= "100000";
            when "1110000111000" => rgb <= "100000";
            when "1110000111001" => rgb <= "100000";
            when "1110000111010" => rgb <= "100000";
            when "1110000111011" => rgb <= "100000";
            when "1110000111100" => rgb <= "100000";
            when "1110000111101" => rgb <= "100000";
            when "1110000111110" => rgb <= "100000";
            when "1110000111111" => rgb <= "100000";
            when "1110001000000" => rgb <= "100000";
            when "1110001000001" => rgb <= "100000";
            when "1110001000010" => rgb <= "100000";
            when "1110001000011" => rgb <= "100000";
            when "1110001000100" => rgb <= "100000";
            when "1110010011100" => rgb <= "010000";
            when "1110010011101" => rgb <= "010000";
            when "1110010011110" => rgb <= "010000";
            when "1110010011111" => rgb <= "010000";
            when "1110010111010" => rgb <= "100000";
            when "1110010111011" => rgb <= "100000";
            when "1110010111100" => rgb <= "100000";
            when "1110010111101" => rgb <= "100000";
            when "1110010111110" => rgb <= "100000";
            when "1110010111111" => rgb <= "100000";
            when "1110011000000" => rgb <= "100000";
            when "1110011000010" => rgb <= "100000";
                    when others => rgb <= "111111";
					-- Don't forget the "others" case!
		end case;
	end if;
end process;
end;


