library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity seven is
  port(
		clk : in std_logic;
		y_in : in  unsigned(5 downto 0);
		x_in : in unsigned(4 downto 0);
		rgb : out std_logic_vector(5 downto 0)
  );
end;
architecture synth of seven is

signal address: std_logic_vector(10 downto 0);

begin
		
address <= std_logic_vector(y_in) & std_logic_vector(x_in);

process (clk)
begin
	if rising_edge(clk) then
			case address is
		            when "00101000001" => rgb <= "001010";
            when "00101000010" => rgb <= "000000";
            when "00101000011" => rgb <= "000000";
            when "00101000100" => rgb <= "000000";
            when "00101000101" => rgb <= "000000";
            when "00101000110" => rgb <= "000000";
            when "00101000111" => rgb <= "000000";
            when "00101001000" => rgb <= "000000";
            when "00101001001" => rgb <= "000000";
            when "00101001010" => rgb <= "000000";
            when "00101001011" => rgb <= "000000";
            when "00101001100" => rgb <= "000000";
            when "00101001101" => rgb <= "000000";
            when "00101001110" => rgb <= "100000";
            when "00101100001" => rgb <= "001010";
            when "00101100010" => rgb <= "000000";
            when "00101100011" => rgb <= "000000";
            when "00101100100" => rgb <= "000000";
            when "00101100101" => rgb <= "000000";
            when "00101100110" => rgb <= "000000";
            when "00101100111" => rgb <= "000000";
            when "00101101000" => rgb <= "000000";
            when "00101101001" => rgb <= "000000";
            when "00101101010" => rgb <= "000000";
            when "00101101011" => rgb <= "000000";
            when "00101101100" => rgb <= "000000";
            when "00101101101" => rgb <= "000000";
            when "00101101110" => rgb <= "100000";
            when "00110000001" => rgb <= "001010";
            when "00110000010" => rgb <= "000000";
            when "00110000011" => rgb <= "000000";
            when "00110000100" => rgb <= "000000";
            when "00110000101" => rgb <= "000000";
            when "00110000110" => rgb <= "000000";
            when "00110000111" => rgb <= "000000";
            when "00110001000" => rgb <= "000000";
            when "00110001001" => rgb <= "000000";
            when "00110001010" => rgb <= "000000";
            when "00110001011" => rgb <= "000000";
            when "00110001100" => rgb <= "000000";
            when "00110001101" => rgb <= "000000";
            when "00110001110" => rgb <= "100000";
            when "00110100001" => rgb <= "001010";
            when "00110100010" => rgb <= "000000";
            when "00110100011" => rgb <= "000000";
            when "00110100100" => rgb <= "000000";
            when "00110100101" => rgb <= "000000";
            when "00110100110" => rgb <= "000000";
            when "00110100111" => rgb <= "000000";
            when "00110101000" => rgb <= "000000";
            when "00110101001" => rgb <= "000000";
            when "00110101010" => rgb <= "000000";
            when "00110101011" => rgb <= "000000";
            when "00110101100" => rgb <= "000000";
            when "00110101101" => rgb <= "000000";
            when "00110101110" => rgb <= "100000";
            when "00111001101" => rgb <= "001010";
            when "00111001110" => rgb <= "000000";
            when "00111001111" => rgb <= "000000";
            when "00111010000" => rgb <= "000000";
            when "00111010001" => rgb <= "000000";
            when "00111010010" => rgb <= "100000";
            when "00111101101" => rgb <= "001010";
            when "00111101110" => rgb <= "000000";
            when "00111101111" => rgb <= "000000";
            when "00111110000" => rgb <= "000000";
            when "00111110001" => rgb <= "000000";
            when "00111110010" => rgb <= "100000";
            when "01000001101" => rgb <= "001010";
            when "01000001110" => rgb <= "000000";
            when "01000001111" => rgb <= "000000";
            when "01000010000" => rgb <= "000000";
            when "01000010001" => rgb <= "000000";
            when "01000010010" => rgb <= "100000";
            when "01000101101" => rgb <= "001010";
            when "01000101110" => rgb <= "000000";
            when "01000101111" => rgb <= "000000";
            when "01000110000" => rgb <= "000000";
            when "01000110001" => rgb <= "000000";
            when "01000110010" => rgb <= "100000";
            when "01001001101" => rgb <= "001010";
            when "01001001110" => rgb <= "000000";
            when "01001001111" => rgb <= "000000";
            when "01001010000" => rgb <= "000000";
            when "01001010001" => rgb <= "000000";
            when "01001010010" => rgb <= "100000";
            when "01001101101" => rgb <= "001010";
            when "01001101110" => rgb <= "000000";
            when "01001101111" => rgb <= "000000";
            when "01001110000" => rgb <= "000000";
            when "01001110001" => rgb <= "000000";
            when "01001110010" => rgb <= "100000";
            when "01010001101" => rgb <= "001010";
            when "01010001110" => rgb <= "000000";
            when "01010001111" => rgb <= "000000";
            when "01010010000" => rgb <= "000000";
            when "01010010001" => rgb <= "000000";
            when "01010010010" => rgb <= "100000";
            when "01010101101" => rgb <= "001010";
            when "01010101110" => rgb <= "000000";
            when "01010101111" => rgb <= "000000";
            when "01010110000" => rgb <= "000000";
            when "01010110001" => rgb <= "000000";
            when "01010110010" => rgb <= "100000";
            when "01011001001" => rgb <= "001010";
            when "01011001010" => rgb <= "000000";
            when "01011001011" => rgb <= "000000";
            when "01011001100" => rgb <= "000000";
            when "01011001101" => rgb <= "000000";
            when "01011001110" => rgb <= "100000";
            when "01011101001" => rgb <= "001010";
            when "01011101010" => rgb <= "000000";
            when "01011101011" => rgb <= "000000";
            when "01011101100" => rgb <= "000000";
            when "01011101101" => rgb <= "000000";
            when "01011101110" => rgb <= "100000";
            when "01100001001" => rgb <= "001010";
            when "01100001010" => rgb <= "000000";
            when "01100001011" => rgb <= "000000";
            when "01100001100" => rgb <= "000000";
            when "01100001101" => rgb <= "000000";
            when "01100001110" => rgb <= "100000";
            when "01100101001" => rgb <= "001010";
            when "01100101010" => rgb <= "000000";
            when "01100101011" => rgb <= "000000";
            when "01100101100" => rgb <= "000000";
            when "01100101101" => rgb <= "000000";
            when "01100101110" => rgb <= "100000";
            when "01101001001" => rgb <= "001010";
            when "01101001010" => rgb <= "000000";
            when "01101001011" => rgb <= "000000";
            when "01101001100" => rgb <= "000000";
            when "01101001101" => rgb <= "000000";
            when "01101001110" => rgb <= "100000";
            when "01101101001" => rgb <= "001010";
            when "01101101010" => rgb <= "000000";
            when "01101101011" => rgb <= "000000";
            when "01101101100" => rgb <= "000000";
            when "01101101101" => rgb <= "000000";
            when "01101101110" => rgb <= "100000";
            when "01110001001" => rgb <= "001010";
            when "01110001010" => rgb <= "000000";
            when "01110001011" => rgb <= "000000";
            when "01110001100" => rgb <= "000000";
            when "01110001101" => rgb <= "000000";
            when "01110001110" => rgb <= "100000";
            when "01110101001" => rgb <= "001010";
            when "01110101010" => rgb <= "000000";
            when "01110101011" => rgb <= "000000";
            when "01110101100" => rgb <= "000000";
            when "01110101101" => rgb <= "000000";
            when "01110101110" => rgb <= "100000";
                    when others => rgb <= "111111";
		end case;
	end if;
end process;
end;